`ifndef CSR__SVH
`define CSR__SVH

`include "isa.svh"

`define CSR__NUM  4096
`define CSR__ALEN $clog2(`CSR__NUM)

`define CSR__RW_FIELD(addr)    addr[11:10]
`define CSR__DEBUG_FIELD(addr) addr[11:4]

`define CSR__READ_ONLY  2'b11
`define CSR__DEBUG_ONLY 8'h7B

`define CSR__CYCLE          12'hC00
`define CSR__CYCLEH         12'hC80
`define CSR__TIME           12'hC01
`define CSR__TIMEH          12'hC81
`define CSR__INSTRET        12'hC02
`define CSR__INSTRETH       12'hC82
`define CSR__HPMCOUNTER3    12'hC03
`define CSR__HPMCOUNTER4    12'hC04
`define CSR__HPMCOUNTER5    12'hC05
`define CSR__HPMCOUNTER6    12'hC06
`define CSR__HPMCOUNTER7    12'hC07
`define CSR__HPMCOUNTER8    12'hC08
`define CSR__HPMCOUNTER9    12'hC09
`define CSR__HPMCOUNTER10   12'hC0A
`define CSR__HPMCOUNTER11   12'hC0B
`define CSR__HPMCOUNTER12   12'hC0C
`define CSR__HPMCOUNTER13   12'hC0D
`define CSR__HPMCOUNTER14   12'hC0E
`define CSR__HPMCOUNTER15   12'hC0F
`define CSR__HPMCOUNTER16   12'hC10
`define CSR__HPMCOUNTER17   12'hC11
`define CSR__HPMCOUNTER18   12'hC12
`define CSR__HPMCOUNTER19   12'hC13
`define CSR__HPMCOUNTER20   12'hC14
`define CSR__HPMCOUNTER21   12'hC15
`define CSR__HPMCOUNTER22   12'hC16
`define CSR__HPMCOUNTER23   12'hC17
`define CSR__HPMCOUNTER24   12'hC18
`define CSR__HPMCOUNTER25   12'hC19
`define CSR__HPMCOUNTER26   12'hC1A
`define CSR__HPMCOUNTER27   12'hC1B
`define CSR__HPMCOUNTER28   12'hC1C
`define CSR__HPMCOUNTER29   12'hC1D
`define CSR__HPMCOUNTER30   12'hC1E
`define CSR__HPMCOUNTER31   12'hC1F
`define CSR__HPMCOUNTER3H   12'hC83
`define CSR__HPMCOUNTER4H   12'hC84
`define CSR__HPMCOUNTER5H   12'hC85
`define CSR__HPMCOUNTER6H   12'hC86
`define CSR__HPMCOUNTER7H   12'hC87
`define CSR__HPMCOUNTER8H   12'hC88
`define CSR__HPMCOUNTER9H   12'hC89
`define CSR__HPMCOUNTER10H  12'hC8A
`define CSR__HPMCOUNTER11H  12'hC8B
`define CSR__HPMCOUNTER12H  12'hC8C
`define CSR__HPMCOUNTER13H  12'hC8D
`define CSR__HPMCOUNTER14H  12'hC8E
`define CSR__HPMCOUNTER15H  12'hC8F
`define CSR__HPMCOUNTER16H  12'hC90
`define CSR__HPMCOUNTER17H  12'hC91
`define CSR__HPMCOUNTER18H  12'hC92
`define CSR__HPMCOUNTER19H  12'hC93
`define CSR__HPMCOUNTER20H  12'hC94
`define CSR__HPMCOUNTER21H  12'hC95
`define CSR__HPMCOUNTER22H  12'hC96
`define CSR__HPMCOUNTER23H  12'hC97
`define CSR__HPMCOUNTER24H  12'hC98
`define CSR__HPMCOUNTER25H  12'hC99
`define CSR__HPMCOUNTER26H  12'hC9A
`define CSR__HPMCOUNTER27H  12'hC9B
`define CSR__HPMCOUNTER28H  12'hC9C
`define CSR__HPMCOUNTER29H  12'hC9D
`define CSR__HPMCOUNTER30H  12'hC9E
`define CSR__HPMCOUNTER31H  12'hC9F
`define CSR__MVENDORID      12'hF11
`define CSR__MARCHID        12'hF12
`define CSR__MIMPID         12'hF13
`define CSR__MHARTID        12'hF14
`define CSR__MCONFIGPTR     12'hF15
`define CSR__MSTATUS        12'h300
`define CSR__MSTATUSH       12'h310
`define CSR__MISA           12'h301
`define CSR__MIE            12'h304
`define CSR__MTVEC          12'h305
`define CSR__MSCRATCH       12'h340
`define CSR__MEPC           12'h341
`define CSR__MCAUSE         12'h342
`define CSR__MTVAL          12'h343
`define CSR__MIP            12'h344
`define CSR__MCYCLE         12'hB00
`define CSR__MCYCLEH        12'hB80
`define CSR__MINSTRET       12'hB02
`define CSR__MINSTRETH      12'hB82
`define CSR__MHPMCOUNTER3   12'hB03
`define CSR__MHPMCOUNTER4   12'hB04
`define CSR__MHPMCOUNTER5   12'hB05
`define CSR__MHPMCOUNTER6   12'hB06
`define CSR__MHPMCOUNTER7   12'hB07
`define CSR__MHPMCOUNTER8   12'hB08
`define CSR__MHPMCOUNTER9   12'hB09
`define CSR__MHPMCOUNTER10  12'hB0A
`define CSR__MHPMCOUNTER11  12'hB0B
`define CSR__MHPMCOUNTER12  12'hB0C
`define CSR__MHPMCOUNTER13  12'hB0D
`define CSR__MHPMCOUNTER14  12'hB0E
`define CSR__MHPMCOUNTER15  12'hB0F
`define CSR__MHPMCOUNTER16  12'hB10
`define CSR__MHPMCOUNTER17  12'hB11
`define CSR__MHPMCOUNTER18  12'hB12
`define CSR__MHPMCOUNTER19  12'hB13
`define CSR__MHPMCOUNTER20  12'hB14
`define CSR__MHPMCOUNTER21  12'hB15
`define CSR__MHPMCOUNTER22  12'hB16
`define CSR__MHPMCOUNTER23  12'hB17
`define CSR__MHPMCOUNTER24  12'hB18
`define CSR__MHPMCOUNTER25  12'hB19
`define CSR__MHPMCOUNTER26  12'hB1A
`define CSR__MHPMCOUNTER27  12'hB1B
`define CSR__MHPMCOUNTER28  12'hB1C
`define CSR__MHPMCOUNTER29  12'hB1D
`define CSR__MHPMCOUNTER30  12'hB1E
`define CSR__MHPMCOUNTER31  12'hB1F
`define CSR__MHPMCOUNTER3H  12'hB83
`define CSR__MHPMCOUNTER4H  12'hB84
`define CSR__MHPMCOUNTER5H  12'hB85
`define CSR__MHPMCOUNTER6H  12'hB86
`define CSR__MHPMCOUNTER7H  12'hB87
`define CSR__MHPMCOUNTER8H  12'hB88
`define CSR__MHPMCOUNTER9H  12'hB89
`define CSR__MHPMCOUNTER10H 12'hB8A
`define CSR__MHPMCOUNTER11H 12'hB8B
`define CSR__MHPMCOUNTER12H 12'hB8C
`define CSR__MHPMCOUNTER13H 12'hB8D
`define CSR__MHPMCOUNTER14H 12'hB8E
`define CSR__MHPMCOUNTER15H 12'hB8F
`define CSR__MHPMCOUNTER16H 12'hB90
`define CSR__MHPMCOUNTER17H 12'hB91
`define CSR__MHPMCOUNTER18H 12'hB92
`define CSR__MHPMCOUNTER19H 12'hB93
`define CSR__MHPMCOUNTER20H 12'hB94
`define CSR__MHPMCOUNTER21H 12'hB95
`define CSR__MHPMCOUNTER22H 12'hB96
`define CSR__MHPMCOUNTER23H 12'hB97
`define CSR__MHPMCOUNTER24H 12'hB98
`define CSR__MHPMCOUNTER25H 12'hB99
`define CSR__MHPMCOUNTER26H 12'hB9A
`define CSR__MHPMCOUNTER27H 12'hB9B
`define CSR__MHPMCOUNTER28H 12'hB9C
`define CSR__MHPMCOUNTER29H 12'hB9D
`define CSR__MHPMCOUNTER30H 12'hB9E
`define CSR__MHPMCOUNTER31H 12'hB9F
`define CSR__MCOUNTINHIBIT  12'h320
`define CSR__MHPMEVENT3     12'h323
`define CSR__MHPMEVENT4     12'h324
`define CSR__MHPMEVENT5     12'h325
`define CSR__MHPMEVENT6     12'h326
`define CSR__MHPMEVENT7     12'h327
`define CSR__MHPMEVENT8     12'h328
`define CSR__MHPMEVENT9     12'h329
`define CSR__MHPMEVENT10    12'h32A
`define CSR__MHPMEVENT11    12'h32B
`define CSR__MHPMEVENT12    12'h32C
`define CSR__MHPMEVENT13    12'h32D
`define CSR__MHPMEVENT14    12'h32E
`define CSR__MHPMEVENT15    12'h32F
`define CSR__MHPMEVENT16    12'h330
`define CSR__MHPMEVENT17    12'h331
`define CSR__MHPMEVENT18    12'h332
`define CSR__MHPMEVENT19    12'h333
`define CSR__MHPMEVENT20    12'h334
`define CSR__MHPMEVENT21    12'h335
`define CSR__MHPMEVENT22    12'h336
`define CSR__MHPMEVENT23    12'h337
`define CSR__MHPMEVENT24    12'h338
`define CSR__MHPMEVENT25    12'h339
`define CSR__MHPMEVENT26    12'h33A
`define CSR__MHPMEVENT27    12'h33B
`define CSR__MHPMEVENT28    12'h33C
`define CSR__MHPMEVENT29    12'h33D
`define CSR__MHPMEVENT30    12'h33E
`define CSR__MHPMEVENT31    12'h33F

`define CSR__WPRI_MASK                 1'b0

`define CSR__CYCLE_MASK               32'h00000000
`define CSR__CYCLEH_MASK              32'h00000000
`define CSR__TIME_MASK                32'h00000000
`define CSR__TIMEH_MASK               32'h00000000
`define CSR__INSTRET_MASK             32'h00000000
`define CSR__INSTRETH_MASK            32'h00000000
`define CSR__HPMCOUNTER3_MASK         32'h00000000
`define CSR__HPMCOUNTER4_MASK         32'h00000000
`define CSR__HPMCOUNTER5_MASK         32'h00000000
`define CSR__HPMCOUNTER6_MASK         32'h00000000
`define CSR__HPMCOUNTER7_MASK         32'h00000000
`define CSR__HPMCOUNTER8_MASK         32'h00000000
`define CSR__HPMCOUNTER9_MASK         32'h00000000
`define CSR__HPMCOUNTER10_MASK        32'h00000000
`define CSR__HPMCOUNTER11_MASK        32'h00000000
`define CSR__HPMCOUNTER12_MASK        32'h00000000
`define CSR__HPMCOUNTER13_MASK        32'h00000000
`define CSR__HPMCOUNTER14_MASK        32'h00000000
`define CSR__HPMCOUNTER15_MASK        32'h00000000
`define CSR__HPMCOUNTER16_MASK        32'h00000000
`define CSR__HPMCOUNTER17_MASK        32'h00000000
`define CSR__HPMCOUNTER18_MASK        32'h00000000
`define CSR__HPMCOUNTER19_MASK        32'h00000000
`define CSR__HPMCOUNTER20_MASK        32'h00000000
`define CSR__HPMCOUNTER21_MASK        32'h00000000
`define CSR__HPMCOUNTER22_MASK        32'h00000000
`define CSR__HPMCOUNTER23_MASK        32'h00000000
`define CSR__HPMCOUNTER24_MASK        32'h00000000
`define CSR__HPMCOUNTER25_MASK        32'h00000000
`define CSR__HPMCOUNTER26_MASK        32'h00000000
`define CSR__HPMCOUNTER27_MASK        32'h00000000
`define CSR__HPMCOUNTER28_MASK        32'h00000000
`define CSR__HPMCOUNTER29_MASK        32'h00000000
`define CSR__HPMCOUNTER30_MASK        32'h00000000
`define CSR__HPMCOUNTER31_MASK        32'h00000000
`define CSR__HPMCOUNTER3H_MASK        32'h00000000
`define CSR__HPMCOUNTER4H_MASK        32'h00000000
`define CSR__HPMCOUNTER5H_MASK        32'h00000000
`define CSR__HPMCOUNTER6H_MASK        32'h00000000
`define CSR__HPMCOUNTER7H_MASK        32'h00000000
`define CSR__HPMCOUNTER8H_MASK        32'h00000000
`define CSR__HPMCOUNTER9H_MASK        32'h00000000
`define CSR__HPMCOUNTER10H_MASK       32'h00000000
`define CSR__HPMCOUNTER11H_MASK       32'h00000000
`define CSR__HPMCOUNTER12H_MASK       32'h00000000
`define CSR__HPMCOUNTER13H_MASK       32'h00000000
`define CSR__HPMCOUNTER14H_MASK       32'h00000000
`define CSR__HPMCOUNTER15H_MASK       32'h00000000
`define CSR__HPMCOUNTER16H_MASK       32'h00000000
`define CSR__HPMCOUNTER17H_MASK       32'h00000000
`define CSR__HPMCOUNTER18H_MASK       32'h00000000
`define CSR__HPMCOUNTER19H_MASK       32'h00000000
`define CSR__HPMCOUNTER20H_MASK       32'h00000000
`define CSR__HPMCOUNTER21H_MASK       32'h00000000
`define CSR__HPMCOUNTER22H_MASK       32'h00000000
`define CSR__HPMCOUNTER23H_MASK       32'h00000000
`define CSR__HPMCOUNTER24H_MASK       32'h00000000
`define CSR__HPMCOUNTER25H_MASK       32'h00000000
`define CSR__HPMCOUNTER26H_MASK       32'h00000000
`define CSR__HPMCOUNTER27H_MASK       32'h00000000
`define CSR__HPMCOUNTER28H_MASK       32'h00000000
`define CSR__HPMCOUNTER29H_MASK       32'h00000000
`define CSR__HPMCOUNTER30H_MASK       32'h00000000
`define CSR__HPMCOUNTER31H_MASK       32'h00000000
`define CSR__MVENDORID_MASK           32'h00000000
`define CSR__MARCHID_MASK             32'h00000000
`define CSR__MIMPID_MASK              32'h00000000
`define CSR__MHARTID_MASK             32'h00000000
`define CSR__MCONFIGPTR_MASK          32'h00000000
`define CSR__MSTATUS_MASK             {`CSR__MSTATUS_SD_MASK,{8{`CSR__WPRI_MASK}},`CSR__MSTATUS_TSR_MASK,`CSR__MSTATUS_TW_MASK,`CSR__MSTATUS_TVM_MASK,`CSR__MSTATUS_MXR_MASK,`CSR__MSTATUS_SUM_MASK,`CSR__MSTATUS_MPRV_MASK,`CSR__MSTATUS_XS_MASK,`CSR__MSTATUS_FS_MASK,`CSR__MSTATUS_MPP_MASK,`CSR__MSTATUS_VS_MASK,`CSR__MSTATUS_SPP_MASK,`CSR__MSTATUS_MPIE_MASK,`CSR__MSTATUS_UBE_MASK,`CSR__MSTATUS_SPIE_MASK,`CSR__WPRI_MASK,`CSR__MSTATUS_MIE_MASK,`CSR__WPRI_MASK,`CSR__MSTATUS_SIE_MASK,`CSR__WPRI_MASK}
`define CSR__MSTATUSH_MASK            {{26{`CSR__WPRI_MASK}},`CSR__MSTATUSH_MBE_MASK,`CSR__MSTATUSH_SBE_MASK,{4{`CSR__WPRI_MASK}}}
`define CSR__MISA_MASK                {`CSR__MISA_MXL_MASK,4'h0,`CSR__MISA_Z_MASK,`CSR__MISA_Y_MASK,`CSR__MISA_X_MASK,`CSR__MISA_W_MASK,`CSR__MISA_V_MASK,`CSR__MISA_U_MASK,`CSR__MISA_T_MASK,`CSR__MISA_S_MASK,`CSR__MISA_R_MASK,`CSR__MISA_Q_MASK,`CSR__MISA_P_MASK,`CSR__MISA_O_MASK,`CSR__MISA_N_MASK,`CSR__MISA_M_MASK,`CSR__MISA_L_MASK,`CSR__MISA_K_MASK,`CSR__MISA_J_MASK,`CSR__MISA_I_MASK,`CSR__MISA_H_MASK,`CSR__MISA_G_MASK,`CSR__MISA_F_MASK,`CSR__MISA_E_MASK,`CSR__MISA_D_MASK,`CSR__MISA_C_MASK,`CSR__MISA_B_MASK,`CSR__MISA_A_MASK}
`define CSR__MIE_MASK                 {16'h0000,4'h0,`CSR__MIE_MEIE_MASK,1'b0,`CSR__MIE_SEIE_MASK,1'b0,`CSR__MIE_MTIE_MASK,1'b0,`CSR__MIE_STIE_MASK,1'b0,`CSR__MIE_MSIE_MASK,1'b0,`CSR__MIE_SSIE_MASK,1'b0}
`define CSR__MTVEC_MASK               {`CSR__MTVEC_BASE_MASK,`CSR__MTVEC_MODE_MASK}
`define CSR__MSCRATCH_MASK            32'hFFFFFFFF
`define CSR__MEPC_MASK                32'hFFFFFFFC
`define CSR__MCAUSE_MASK              {`CSR__MCAUSE_INT_MASK,`CSR__MCAUSE_CODE_MASK}
`define CSR__MTVAL_MASK               32'hFFFFFFFF
`define CSR__MIP_MASK                 {16'h0000,4'h0,`CSR__MIP_MEIP_MASK,1'b0,`CSR__MIP_SEIP_MASK,1'b0,`CSR__MIP_MTIP_MASK,1'b0,`CSR__MIP_STIP_MASK,1'b0,`CSR__MIP_MSIP_MASK,1'b0,`CSR__MIP_SSIP_MASK,1'b0}
`define CSR__MCYCLE_MASK              32'hFFFFFFFF
`define CSR__MCYCLEH_MASK             32'hFFFFFFFF
`define CSR__MINSTRET_MASK            32'hFFFFFFFF
`define CSR__MINSTRETH_MASK           32'hFFFFFFFF
`define CSR__MHPMCOUNTER3_MASK        32'h00000000
`define CSR__MHPMCOUNTER4_MASK        32'h00000000
`define CSR__MHPMCOUNTER5_MASK        32'h00000000
`define CSR__MHPMCOUNTER6_MASK        32'h00000000
`define CSR__MHPMCOUNTER7_MASK        32'h00000000
`define CSR__MHPMCOUNTER8_MASK        32'h00000000
`define CSR__MHPMCOUNTER9_MASK        32'h00000000
`define CSR__MHPMCOUNTER10_MASK       32'h00000000
`define CSR__MHPMCOUNTER11_MASK       32'h00000000
`define CSR__MHPMCOUNTER12_MASK       32'h00000000
`define CSR__MHPMCOUNTER13_MASK       32'h00000000
`define CSR__MHPMCOUNTER14_MASK       32'h00000000
`define CSR__MHPMCOUNTER15_MASK       32'h00000000
`define CSR__MHPMCOUNTER16_MASK       32'h00000000
`define CSR__MHPMCOUNTER17_MASK       32'h00000000
`define CSR__MHPMCOUNTER18_MASK       32'h00000000
`define CSR__MHPMCOUNTER19_MASK       32'h00000000
`define CSR__MHPMCOUNTER20_MASK       32'h00000000
`define CSR__MHPMCOUNTER21_MASK       32'h00000000
`define CSR__MHPMCOUNTER22_MASK       32'h00000000
`define CSR__MHPMCOUNTER23_MASK       32'h00000000
`define CSR__MHPMCOUNTER24_MASK       32'h00000000
`define CSR__MHPMCOUNTER25_MASK       32'h00000000
`define CSR__MHPMCOUNTER26_MASK       32'h00000000
`define CSR__MHPMCOUNTER27_MASK       32'h00000000
`define CSR__MHPMCOUNTER28_MASK       32'h00000000
`define CSR__MHPMCOUNTER29_MASK       32'h00000000
`define CSR__MHPMCOUNTER30_MASK       32'h00000000
`define CSR__MHPMCOUNTER31_MASK       32'h00000000
`define CSR__MHPMCOUNTER3H_MASK       32'h00000000
`define CSR__MHPMCOUNTER4H_MASK       32'h00000000
`define CSR__MHPMCOUNTER5H_MASK       32'h00000000
`define CSR__MHPMCOUNTER6H_MASK       32'h00000000
`define CSR__MHPMCOUNTER7H_MASK       32'h00000000
`define CSR__MHPMCOUNTER8H_MASK       32'h00000000
`define CSR__MHPMCOUNTER9H_MASK       32'h00000000
`define CSR__MHPMCOUNTER10H_MASK      32'h00000000
`define CSR__MHPMCOUNTER11H_MASK      32'h00000000
`define CSR__MHPMCOUNTER12H_MASK      32'h00000000
`define CSR__MHPMCOUNTER13H_MASK      32'h00000000
`define CSR__MHPMCOUNTER14H_MASK      32'h00000000
`define CSR__MHPMCOUNTER15H_MASK      32'h00000000
`define CSR__MHPMCOUNTER16H_MASK      32'h00000000
`define CSR__MHPMCOUNTER17H_MASK      32'h00000000
`define CSR__MHPMCOUNTER18H_MASK      32'h00000000
`define CSR__MHPMCOUNTER19H_MASK      32'h00000000
`define CSR__MHPMCOUNTER20H_MASK      32'h00000000
`define CSR__MHPMCOUNTER21H_MASK      32'h00000000
`define CSR__MHPMCOUNTER22H_MASK      32'h00000000
`define CSR__MHPMCOUNTER23H_MASK      32'h00000000
`define CSR__MHPMCOUNTER24H_MASK      32'h00000000
`define CSR__MHPMCOUNTER25H_MASK      32'h00000000
`define CSR__MHPMCOUNTER26H_MASK      32'h00000000
`define CSR__MHPMCOUNTER27H_MASK      32'h00000000
`define CSR__MHPMCOUNTER28H_MASK      32'h00000000
`define CSR__MHPMCOUNTER29H_MASK      32'h00000000
`define CSR__MHPMCOUNTER30H_MASK      32'h00000000
`define CSR__MHPMCOUNTER31H_MASK      32'h00000000
`define CSR__MCOUNTINHIBIT_MASK       {`CSR__MCOUNTINHIBIT_HPM31_MASK,`CSR__MCOUNTINHIBIT_HPM30_MASK,`CSR__MCOUNTINHIBIT_HPM29_MASK,`CSR__MCOUNTINHIBIT_HPM28_MASK,`CSR__MCOUNTINHIBIT_HPM27_MASK,`CSR__MCOUNTINHIBIT_HPM26_MASK,`CSR__MCOUNTINHIBIT_HPM25_MASK,`CSR__MCOUNTINHIBIT_HPM24_MASK,`CSR__MCOUNTINHIBIT_HPM23_MASK,`CSR__MCOUNTINHIBIT_HPM22_MASK,`CSR__MCOUNTINHIBIT_HPM21_MASK,`CSR__MCOUNTINHIBIT_HPM20_MASK,`CSR__MCOUNTINHIBIT_HPM19_MASK,`CSR__MCOUNTINHIBIT_HPM18_MASK,`CSR__MCOUNTINHIBIT_HPM17_MASK,`CSR__MCOUNTINHIBIT_HPM16_MASK,`CSR__MCOUNTINHIBIT_HPM15_MASK,`CSR__MCOUNTINHIBIT_HPM14_MASK,`CSR__MCOUNTINHIBIT_HPM13_MASK,`CSR__MCOUNTINHIBIT_HPM12_MASK,`CSR__MCOUNTINHIBIT_HPM11_MASK,`CSR__MCOUNTINHIBIT_HPM10_MASK,`CSR__MCOUNTINHIBIT_HPM9_MASK,`CSR__MCOUNTINHIBIT_HPM8_MASK,`CSR__MCOUNTINHIBIT_HPM7_MASK,`CSR__MCOUNTINHIBIT_HPM6_MASK,`CSR__MCOUNTINHIBIT_HPM5_MASK,`CSR__MCOUNTINHIBIT_HPM4_MASK,`CSR__MCOUNTINHIBIT_HPM3_MASK,`CSR__MCOUNTINHIBIT_IR_MASK,1'b0,`CSR__MCOUNTINHIBIT_CY_MASK}
`define CSR__MHPMEVENT3_MASK          32'h00000000
`define CSR__MHPMEVENT4_MASK          32'h00000000
`define CSR__MHPMEVENT5_MASK          32'h00000000
`define CSR__MHPMEVENT6_MASK          32'h00000000
`define CSR__MHPMEVENT7_MASK          32'h00000000
`define CSR__MHPMEVENT8_MASK          32'h00000000
`define CSR__MHPMEVENT9_MASK          32'h00000000
`define CSR__MHPMEVENT10_MASK         32'h00000000
`define CSR__MHPMEVENT11_MASK         32'h00000000
`define CSR__MHPMEVENT12_MASK         32'h00000000
`define CSR__MHPMEVENT13_MASK         32'h00000000
`define CSR__MHPMEVENT14_MASK         32'h00000000
`define CSR__MHPMEVENT15_MASK         32'h00000000
`define CSR__MHPMEVENT16_MASK         32'h00000000
`define CSR__MHPMEVENT17_MASK         32'h00000000
`define CSR__MHPMEVENT18_MASK         32'h00000000
`define CSR__MHPMEVENT19_MASK         32'h00000000
`define CSR__MHPMEVENT20_MASK         32'h00000000
`define CSR__MHPMEVENT21_MASK         32'h00000000
`define CSR__MHPMEVENT22_MASK         32'h00000000
`define CSR__MHPMEVENT23_MASK         32'h00000000
`define CSR__MHPMEVENT24_MASK         32'h00000000
`define CSR__MHPMEVENT25_MASK         32'h00000000
`define CSR__MHPMEVENT26_MASK         32'h00000000
`define CSR__MHPMEVENT27_MASK         32'h00000000
`define CSR__MHPMEVENT28_MASK         32'h00000000
`define CSR__MHPMEVENT29_MASK         32'h00000000
`define CSR__MHPMEVENT30_MASK         32'h00000000
`define CSR__MHPMEVENT31_MASK         32'h00000000

`define CSR__MISA_MXL_MASK             2'b00
`define CSR__MISA_A_MASK               1'b0
`define CSR__MISA_B_MASK               1'b0
`define CSR__MISA_C_MASK               1'b0
`define CSR__MISA_D_MASK               1'b0
`define CSR__MISA_E_MASK               1'b0
`define CSR__MISA_F_MASK               1'b0
`define CSR__MISA_G_MASK               1'b0
`define CSR__MISA_H_MASK               1'b0
`define CSR__MISA_I_MASK               1'b0
`define CSR__MISA_J_MASK               1'b0
`define CSR__MISA_K_MASK               1'b0
`define CSR__MISA_L_MASK               1'b0
`define CSR__MISA_M_MASK               1'b0
`define CSR__MISA_N_MASK               1'b0
`define CSR__MISA_O_MASK               1'b0
`define CSR__MISA_P_MASK               1'b0
`define CSR__MISA_Q_MASK               1'b0
`define CSR__MISA_R_MASK               1'b0
`define CSR__MISA_S_MASK               1'b0
`define CSR__MISA_T_MASK               1'b0
`define CSR__MISA_U_MASK               1'b0
`define CSR__MISA_V_MASK               1'b0
`define CSR__MISA_W_MASK               1'b0
`define CSR__MISA_X_MASK               1'b0
`define CSR__MISA_Y_MASK               1'b0
`define CSR__MISA_Z_MASK               1'b0

`define CSR__MSTATUS_SD_MASK           1'b0
`define CSR__MSTATUS_TSR_MASK          1'b0
`define CSR__MSTATUS_TW_MASK           1'b0
`define CSR__MSTATUS_TVM_MASK          1'b0
`define CSR__MSTATUS_MXR_MASK          1'b0
`define CSR__MSTATUS_SUM_MASK          1'b0
`define CSR__MSTATUS_MPRV_MASK         1'b0
`define CSR__MSTATUS_XS_MASK           2'b00
`define CSR__MSTATUS_FS_MASK           2'b00
`define CSR__MSTATUS_MPP_MASK          2'b00
`define CSR__MSTATUS_VS_MASK           2'b00
`define CSR__MSTATUS_SPP_MASK          1'b0
`define CSR__MSTATUS_MPIE_MASK         1'b1
`define CSR__MSTATUS_UBE_MASK          1'b0
`define CSR__MSTATUS_SPIE_MASK         1'b0
`define CSR__MSTATUS_MIE_MASK          1'b1
`define CSR__MSTATUS_SIE_MASK          1'b0

`define CSR__MSTATUSH_MBE_MASK         1'b0
`define CSR__MSTATUSH_SBE_MASK         1'b0

`define CSR__MTVEC_BASE_MASK          30'hFFFFFFFF
`define CSR__MTVEC_MODE_MASK           2'b01

`define CSR__MIP_MEIP_MASK             1'b0
`define CSR__MIP_SEIP_MASK             1'b0
`define CSR__MIP_MTIP_MASK             1'b0
`define CSR__MIP_STIP_MASK             1'b0
`define CSR__MIP_MSIP_MASK             1'b0
`define CSR__MIP_SSIP_MASK             1'b0

`define CSR__MIE_MEIE_MASK             1'b1
`define CSR__MIE_SEIE_MASK             1'b0
`define CSR__MIE_MTIE_MASK             1'b1
`define CSR__MIE_STIE_MASK             1'b0
`define CSR__MIE_MSIE_MASK             1'b0
`define CSR__MIE_SSIE_MASK             1'b0

`define CSR__MCOUNTINHIBIT_CY_MASK     1'b1
`define CSR__MCOUNTINHIBIT_IR_MASK     1'b1
`define CSR__MCOUNTINHIBIT_HPM3_MASK   1'b0
`define CSR__MCOUNTINHIBIT_HPM4_MASK   1'b0
`define CSR__MCOUNTINHIBIT_HPM5_MASK   1'b0
`define CSR__MCOUNTINHIBIT_HPM6_MASK   1'b0
`define CSR__MCOUNTINHIBIT_HPM7_MASK   1'b0
`define CSR__MCOUNTINHIBIT_HPM8_MASK   1'b0
`define CSR__MCOUNTINHIBIT_HPM9_MASK   1'b0
`define CSR__MCOUNTINHIBIT_HPM10_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM11_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM12_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM13_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM14_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM15_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM16_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM17_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM18_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM19_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM20_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM21_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM22_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM23_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM24_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM25_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM26_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM27_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM28_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM29_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM30_MASK  1'b0
`define CSR__MCOUNTINHIBIT_HPM31_MASK  1'b0

`define CSR__MCAUSE_INT_MASK           1'b1
`define CSR__MCAUSE_CODE_MASK         31'hFFFFFFFF

`define CSR__WPRI_VALUE                 1'b0

`define CSR__CYCLE_VALUE               32'h00000000
`define CSR__CYCLEH_VALUE              32'h00000000
`define CSR__TIME_VALUE                32'h00000000
`define CSR__TIMEH_VALUE               32'h00000000
`define CSR__INSTRET_VALUE             32'h00000000
`define CSR__INSTRETH_VALUE            32'h00000000
`define CSR__HPMCOUNTER3_VALUE         32'h00000000
`define CSR__HPMCOUNTER4_VALUE         32'h00000000
`define CSR__HPMCOUNTER5_VALUE         32'h00000000
`define CSR__HPMCOUNTER6_VALUE         32'h00000000
`define CSR__HPMCOUNTER7_VALUE         32'h00000000
`define CSR__HPMCOUNTER8_VALUE         32'h00000000
`define CSR__HPMCOUNTER9_VALUE         32'h00000000
`define CSR__HPMCOUNTER10_VALUE        32'h00000000
`define CSR__HPMCOUNTER11_VALUE        32'h00000000
`define CSR__HPMCOUNTER12_VALUE        32'h00000000
`define CSR__HPMCOUNTER13_VALUE        32'h00000000
`define CSR__HPMCOUNTER14_VALUE        32'h00000000
`define CSR__HPMCOUNTER15_VALUE        32'h00000000
`define CSR__HPMCOUNTER16_VALUE        32'h00000000
`define CSR__HPMCOUNTER17_VALUE        32'h00000000
`define CSR__HPMCOUNTER18_VALUE        32'h00000000
`define CSR__HPMCOUNTER19_VALUE        32'h00000000
`define CSR__HPMCOUNTER20_VALUE        32'h00000000
`define CSR__HPMCOUNTER21_VALUE        32'h00000000
`define CSR__HPMCOUNTER22_VALUE        32'h00000000
`define CSR__HPMCOUNTER23_VALUE        32'h00000000
`define CSR__HPMCOUNTER24_VALUE        32'h00000000
`define CSR__HPMCOUNTER25_VALUE        32'h00000000
`define CSR__HPMCOUNTER26_VALUE        32'h00000000
`define CSR__HPMCOUNTER27_VALUE        32'h00000000
`define CSR__HPMCOUNTER28_VALUE        32'h00000000
`define CSR__HPMCOUNTER29_VALUE        32'h00000000
`define CSR__HPMCOUNTER30_VALUE        32'h00000000
`define CSR__HPMCOUNTER31_VALUE        32'h00000000
`define CSR__HPMCOUNTER3H_VALUE        32'h00000000
`define CSR__HPMCOUNTER4H_VALUE        32'h00000000
`define CSR__HPMCOUNTER5H_VALUE        32'h00000000
`define CSR__HPMCOUNTER6H_VALUE        32'h00000000
`define CSR__HPMCOUNTER7H_VALUE        32'h00000000
`define CSR__HPMCOUNTER8H_VALUE        32'h00000000
`define CSR__HPMCOUNTER9H_VALUE        32'h00000000
`define CSR__HPMCOUNTER10H_VALUE       32'h00000000
`define CSR__HPMCOUNTER11H_VALUE       32'h00000000
`define CSR__HPMCOUNTER12H_VALUE       32'h00000000
`define CSR__HPMCOUNTER13H_VALUE       32'h00000000
`define CSR__HPMCOUNTER14H_VALUE       32'h00000000
`define CSR__HPMCOUNTER15H_VALUE       32'h00000000
`define CSR__HPMCOUNTER16H_VALUE       32'h00000000
`define CSR__HPMCOUNTER17H_VALUE       32'h00000000
`define CSR__HPMCOUNTER18H_VALUE       32'h00000000
`define CSR__HPMCOUNTER19H_VALUE       32'h00000000
`define CSR__HPMCOUNTER20H_VALUE       32'h00000000
`define CSR__HPMCOUNTER21H_VALUE       32'h00000000
`define CSR__HPMCOUNTER22H_VALUE       32'h00000000
`define CSR__HPMCOUNTER23H_VALUE       32'h00000000
`define CSR__HPMCOUNTER24H_VALUE       32'h00000000
`define CSR__HPMCOUNTER25H_VALUE       32'h00000000
`define CSR__HPMCOUNTER26H_VALUE       32'h00000000
`define CSR__HPMCOUNTER27H_VALUE       32'h00000000
`define CSR__HPMCOUNTER28H_VALUE       32'h00000000
`define CSR__HPMCOUNTER29H_VALUE       32'h00000000
`define CSR__HPMCOUNTER30H_VALUE       32'h00000000
`define CSR__HPMCOUNTER31H_VALUE       32'h00000000
`define CSR__MVENDORID_VALUE           32'h00000000
`define CSR__MARCHID_VALUE             32'h00000000
`define CSR__MIMPID_VALUE              32'h00000000
`define CSR__MHARTID_VALUE             32'h00000000
`define CSR__MCONFIGPTR_VALUE          32'h00000000
`define CSR__MSTATUS_VALUE             {`CSR__MSTATUS_SD_VALUE,{8{`CSR__WPRI_VALUE}},`CSR__MSTATUS_TSR_VALUE,`CSR__MSTATUS_TW_VALUE,`CSR__MSTATUS_TVM_VALUE,`CSR__MSTATUS_MXR_VALUE,`CSR__MSTATUS_SUM_VALUE,`CSR__MSTATUS_MPRV_VALUE,`CSR__MSTATUS_XS_VALUE,`CSR__MSTATUS_FS_VALUE,`CSR__MSTATUS_MPP_VALUE,`CSR__MSTATUS_VS_VALUE,`CSR__MSTATUS_SPP_VALUE,`CSR__MSTATUS_MPIE_VALUE,`CSR__MSTATUS_UBE_VALUE,`CSR__MSTATUS_SPIE_VALUE,`CSR__WPRI_VALUE,`CSR__MSTATUS_MIE_VALUE,`CSR__WPRI_VALUE,`CSR__MSTATUS_SIE_VALUE,`CSR__WPRI_VALUE}
`define CSR__MSTATUSH_VALUE            {{26{`CSR__WPRI_VALUE}},`CSR__MSTATUSH_MBE_VALUE,`CSR__MSTATUSH_SBE_VALUE,{4{`CSR__WPRI_VALUE}}}
`define CSR__MISA_VALUE                {`CSR__MISA_MXL_VALUE,4'h0,`CSR__MISA_Z_VALUE,`CSR__MISA_Y_VALUE,`CSR__MISA_X_VALUE,`CSR__MISA_W_VALUE,`CSR__MISA_V_VALUE,`CSR__MISA_U_VALUE,`CSR__MISA_T_VALUE,`CSR__MISA_S_VALUE,`CSR__MISA_R_VALUE,`CSR__MISA_Q_VALUE,`CSR__MISA_P_VALUE,`CSR__MISA_O_VALUE,`CSR__MISA_N_VALUE,`CSR__MISA_M_VALUE,`CSR__MISA_L_VALUE,`CSR__MISA_K_VALUE,`CSR__MISA_J_VALUE,`CSR__MISA_I_VALUE,`CSR__MISA_H_VALUE,`CSR__MISA_G_VALUE,`CSR__MISA_F_VALUE,`CSR__MISA_E_VALUE,`CSR__MISA_D_VALUE,`CSR__MISA_C_VALUE,`CSR__MISA_B_VALUE,`CSR__MISA_A_VALUE}
`define CSR__MIE_VALUE                 {16'h0000,4'h0,`CSR__MIE_MEIE_VALUE,1'b0,`CSR__MIE_SEIE_VALUE,1'b0,`CSR__MIE_MTIE_VALUE,1'b0,`CSR__MIE_STIE_VALUE,1'b0,`CSR__MIE_MSIE_VALUE,1'b0,`CSR__MIE_SSIE_VALUE,1'b0}
`define CSR__MTVEC_VALUE               {`CSR__MTVEC_BASE_VALUE,`CSR__MTVEC_MODE_VALUE}
`define CSR__MSCRATCH_VALUE            32'h00000000
`define CSR__MEPC_VALUE                32'h00000000
`define CSR__MCAUSE_VALUE              {`CSR__MCAUSE_INT_VALUE,`CSR__MCAUSE_CODE_VALUE}
`define CSR__MTVAL_VALUE               32'h00000000
`define CSR__MIP_VALUE                 {16'h0000,4'h0,`CSR__MIP_MEIP_VALUE,1'b0,`CSR__MIP_SEIP_VALUE,1'b0,`CSR__MIP_MTIP_VALUE,1'b0,`CSR__MIP_STIP_VALUE,1'b0,`CSR__MIP_MSIP_VALUE,1'b0,`CSR__MIP_SSIP_VALUE,1'b0}
`define CSR__MCYCLE_VALUE              32'h00000000
`define CSR__MCYCLEH_VALUE             32'h00000000
`define CSR__MINSTRET_VALUE            32'h00000000
`define CSR__MINSTRETH_VALUE           32'h00000000
`define CSR__MHPMCOUNTER3_VALUE        32'h00000000
`define CSR__MHPMCOUNTER4_VALUE        32'h00000000
`define CSR__MHPMCOUNTER5_VALUE        32'h00000000
`define CSR__MHPMCOUNTER6_VALUE        32'h00000000
`define CSR__MHPMCOUNTER7_VALUE        32'h00000000
`define CSR__MHPMCOUNTER8_VALUE        32'h00000000
`define CSR__MHPMCOUNTER9_VALUE        32'h00000000
`define CSR__MHPMCOUNTER10_VALUE       32'h00000000
`define CSR__MHPMCOUNTER11_VALUE       32'h00000000
`define CSR__MHPMCOUNTER12_VALUE       32'h00000000
`define CSR__MHPMCOUNTER13_VALUE       32'h00000000
`define CSR__MHPMCOUNTER14_VALUE       32'h00000000
`define CSR__MHPMCOUNTER15_VALUE       32'h00000000
`define CSR__MHPMCOUNTER16_VALUE       32'h00000000
`define CSR__MHPMCOUNTER17_VALUE       32'h00000000
`define CSR__MHPMCOUNTER18_VALUE       32'h00000000
`define CSR__MHPMCOUNTER19_VALUE       32'h00000000
`define CSR__MHPMCOUNTER20_VALUE       32'h00000000
`define CSR__MHPMCOUNTER21_VALUE       32'h00000000
`define CSR__MHPMCOUNTER22_VALUE       32'h00000000
`define CSR__MHPMCOUNTER23_VALUE       32'h00000000
`define CSR__MHPMCOUNTER24_VALUE       32'h00000000
`define CSR__MHPMCOUNTER25_VALUE       32'h00000000
`define CSR__MHPMCOUNTER26_VALUE       32'h00000000
`define CSR__MHPMCOUNTER27_VALUE       32'h00000000
`define CSR__MHPMCOUNTER28_VALUE       32'h00000000
`define CSR__MHPMCOUNTER29_VALUE       32'h00000000
`define CSR__MHPMCOUNTER30_VALUE       32'h00000000
`define CSR__MHPMCOUNTER31_VALUE       32'h00000000
`define CSR__MHPMCOUNTER3H_VALUE       32'h00000000
`define CSR__MHPMCOUNTER4H_VALUE       32'h00000000
`define CSR__MHPMCOUNTER5H_VALUE       32'h00000000
`define CSR__MHPMCOUNTER6H_VALUE       32'h00000000
`define CSR__MHPMCOUNTER7H_VALUE       32'h00000000
`define CSR__MHPMCOUNTER8H_VALUE       32'h00000000
`define CSR__MHPMCOUNTER9H_VALUE       32'h00000000
`define CSR__MHPMCOUNTER10H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER11H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER12H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER13H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER14H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER15H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER16H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER17H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER18H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER19H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER20H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER21H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER22H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER23H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER24H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER25H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER26H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER27H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER28H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER29H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER30H_VALUE      32'h00000000
`define CSR__MHPMCOUNTER31H_VALUE      32'h00000000
`define CSR__MCOUNTINHIBIT_VALUE       {`CSR__MCOUNTINHIBIT_HPM31_VALUE,`CSR__MCOUNTINHIBIT_HPM30_VALUE,`CSR__MCOUNTINHIBIT_HPM29_VALUE,`CSR__MCOUNTINHIBIT_HPM28_VALUE,`CSR__MCOUNTINHIBIT_HPM27_VALUE,`CSR__MCOUNTINHIBIT_HPM26_VALUE,`CSR__MCOUNTINHIBIT_HPM25_VALUE,`CSR__MCOUNTINHIBIT_HPM24_VALUE,`CSR__MCOUNTINHIBIT_HPM23_VALUE,`CSR__MCOUNTINHIBIT_HPM22_VALUE,`CSR__MCOUNTINHIBIT_HPM21_VALUE,`CSR__MCOUNTINHIBIT_HPM20_VALUE,`CSR__MCOUNTINHIBIT_HPM19_VALUE,`CSR__MCOUNTINHIBIT_HPM18_VALUE,`CSR__MCOUNTINHIBIT_HPM17_VALUE,`CSR__MCOUNTINHIBIT_HPM16_VALUE,`CSR__MCOUNTINHIBIT_HPM15_VALUE,`CSR__MCOUNTINHIBIT_HPM14_VALUE,`CSR__MCOUNTINHIBIT_HPM13_VALUE,`CSR__MCOUNTINHIBIT_HPM12_VALUE,`CSR__MCOUNTINHIBIT_HPM11_VALUE,`CSR__MCOUNTINHIBIT_HPM10_VALUE,`CSR__MCOUNTINHIBIT_HPM9_VALUE,`CSR__MCOUNTINHIBIT_HPM8_VALUE,`CSR__MCOUNTINHIBIT_HPM7_VALUE,`CSR__MCOUNTINHIBIT_HPM6_VALUE,`CSR__MCOUNTINHIBIT_HPM5_VALUE,`CSR__MCOUNTINHIBIT_HPM4_VALUE,`CSR__MCOUNTINHIBIT_HPM3_VALUE,`CSR__MCOUNTINHIBIT_IR_VALUE,1'b0,`CSR__MCOUNTINHIBIT_CY_VALUE}
`define CSR__MHPMEVENT3_VALUE          32'h00000000
`define CSR__MHPMEVENT4_VALUE          32'h00000000
`define CSR__MHPMEVENT5_VALUE          32'h00000000
`define CSR__MHPMEVENT6_VALUE          32'h00000000
`define CSR__MHPMEVENT7_VALUE          32'h00000000
`define CSR__MHPMEVENT8_VALUE          32'h00000000
`define CSR__MHPMEVENT9_VALUE          32'h00000000
`define CSR__MHPMEVENT10_VALUE         32'h00000000
`define CSR__MHPMEVENT11_VALUE         32'h00000000
`define CSR__MHPMEVENT12_VALUE         32'h00000000
`define CSR__MHPMEVENT13_VALUE         32'h00000000
`define CSR__MHPMEVENT14_VALUE         32'h00000000
`define CSR__MHPMEVENT15_VALUE         32'h00000000
`define CSR__MHPMEVENT16_VALUE         32'h00000000
`define CSR__MHPMEVENT17_VALUE         32'h00000000
`define CSR__MHPMEVENT18_VALUE         32'h00000000
`define CSR__MHPMEVENT19_VALUE         32'h00000000
`define CSR__MHPMEVENT20_VALUE         32'h00000000
`define CSR__MHPMEVENT21_VALUE         32'h00000000
`define CSR__MHPMEVENT22_VALUE         32'h00000000
`define CSR__MHPMEVENT23_VALUE         32'h00000000
`define CSR__MHPMEVENT24_VALUE         32'h00000000
`define CSR__MHPMEVENT25_VALUE         32'h00000000
`define CSR__MHPMEVENT26_VALUE         32'h00000000
`define CSR__MHPMEVENT27_VALUE         32'h00000000
`define CSR__MHPMEVENT28_VALUE         32'h00000000
`define CSR__MHPMEVENT29_VALUE         32'h00000000
`define CSR__MHPMEVENT30_VALUE         32'h00000000
`define CSR__MHPMEVENT31_VALUE         32'h00000000

`define CSR__MISA_MXL_VALUE             2'b01
`define CSR__MISA_A_VALUE               1'b0
`define CSR__MISA_B_VALUE               1'b0
`define CSR__MISA_C_VALUE               1'b0
`define CSR__MISA_D_VALUE               1'b0
`define CSR__MISA_E_VALUE               1'b0
`define CSR__MISA_F_VALUE               1'b0
`define CSR__MISA_G_VALUE               1'b0
`define CSR__MISA_H_VALUE               1'b0
`define CSR__MISA_I_VALUE               1'b1
`define CSR__MISA_J_VALUE               1'b0
`define CSR__MISA_K_VALUE               1'b0
`define CSR__MISA_L_VALUE               1'b0
`define CSR__MISA_M_VALUE               `ISA__MEXT
`define CSR__MISA_N_VALUE               1'b0
`define CSR__MISA_O_VALUE               1'b0
`define CSR__MISA_P_VALUE               1'b0
`define CSR__MISA_Q_VALUE               1'b0
`define CSR__MISA_R_VALUE               1'b0
`define CSR__MISA_S_VALUE               1'b0
`define CSR__MISA_T_VALUE               1'b0
`define CSR__MISA_U_VALUE               1'b0
`define CSR__MISA_V_VALUE               1'b0
`define CSR__MISA_W_VALUE               1'b0
`define CSR__MISA_X_VALUE               1'b0
`define CSR__MISA_Y_VALUE               1'b0
`define CSR__MISA_Z_VALUE               1'b0

`define CSR__MSTATUS_SD_VALUE           1'b0
`define CSR__MSTATUS_TSR_VALUE          1'b0
`define CSR__MSTATUS_TW_VALUE           1'b0
`define CSR__MSTATUS_TVM_VALUE          1'b0
`define CSR__MSTATUS_MXR_VALUE          1'b0
`define CSR__MSTATUS_SUM_VALUE          1'b0
`define CSR__MSTATUS_MPRV_VALUE         1'b0
`define CSR__MSTATUS_XS_VALUE           2'b00
`define CSR__MSTATUS_FS_VALUE           2'b00
`define CSR__MSTATUS_MPP_VALUE          2'b11
`define CSR__MSTATUS_VS_VALUE           2'b00
`define CSR__MSTATUS_SPP_VALUE          1'b0
`define CSR__MSTATUS_MPIE_VALUE         1'b0
`define CSR__MSTATUS_UBE_VALUE          1'b0
`define CSR__MSTATUS_SPIE_VALUE         1'b0
`define CSR__MSTATUS_MIE_VALUE          1'b0
`define CSR__MSTATUS_SIE_VALUE          1'b0

`define CSR__MSTATUSH_MBE_VALUE         1'b0
`define CSR__MSTATUSH_SBE_VALUE         1'b0

`define CSR__MTVEC_BASE_VALUE          30'h00000000
`define CSR__MTVEC_MODE_VALUE           2'b00

`define CSR__MIP_MEIP_VALUE             1'b0
`define CSR__MIP_SEIP_VALUE             1'b0
`define CSR__MIP_MTIP_VALUE             1'b0
`define CSR__MIP_STIP_VALUE             1'b0
`define CSR__MIP_MSIP_VALUE             1'b0
`define CSR__MIP_SSIP_VALUE             1'b0

`define CSR__MIE_MEIE_VALUE             1'b0
`define CSR__MIE_SEIE_VALUE             1'b0
`define CSR__MIE_MTIE_VALUE             1'b0
`define CSR__MIE_STIE_VALUE             1'b0
`define CSR__MIE_MSIE_VALUE             1'b0
`define CSR__MIE_SSIE_VALUE             1'b0

`define CSR__MCOUNTINHIBIT_CY_VALUE     1'b0
`define CSR__MCOUNTINHIBIT_IR_VALUE     1'b0
`define CSR__MCOUNTINHIBIT_HPM3_VALUE   1'b0
`define CSR__MCOUNTINHIBIT_HPM4_VALUE   1'b0
`define CSR__MCOUNTINHIBIT_HPM5_VALUE   1'b0
`define CSR__MCOUNTINHIBIT_HPM6_VALUE   1'b0
`define CSR__MCOUNTINHIBIT_HPM7_VALUE   1'b0
`define CSR__MCOUNTINHIBIT_HPM8_VALUE   1'b0
`define CSR__MCOUNTINHIBIT_HPM9_VALUE   1'b0
`define CSR__MCOUNTINHIBIT_HPM10_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM11_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM12_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM13_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM14_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM15_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM16_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM17_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM18_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM19_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM20_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM21_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM22_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM23_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM24_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM25_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM26_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM27_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM28_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM29_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM30_VALUE  1'b0
`define CSR__MCOUNTINHIBIT_HPM31_VALUE  1'b0

`define CSR__MCAUSE_INT_VALUE           1'b0
`define CSR__MCAUSE_CODE_VALUE         31'h00000000



`define CSRGEN__FOREACH(TARGET) \
`TARGET(CYCLE)          \
`TARGET(CYCLEH)         \
`TARGET(TIME)           \
`TARGET(TIMEH)          \
`TARGET(INSTRET)        \
`TARGET(INSTRETH)       \
`TARGET(HPMCOUNTER3)    \
`TARGET(HPMCOUNTER4)    \
`TARGET(HPMCOUNTER5)    \
`TARGET(HPMCOUNTER6)    \
`TARGET(HPMCOUNTER7)    \
`TARGET(HPMCOUNTER8)    \
`TARGET(HPMCOUNTER9)    \
`TARGET(HPMCOUNTER10)   \
`TARGET(HPMCOUNTER11)   \
`TARGET(HPMCOUNTER12)   \
`TARGET(HPMCOUNTER13)   \
`TARGET(HPMCOUNTER14)   \
`TARGET(HPMCOUNTER15)   \
`TARGET(HPMCOUNTER16)   \
`TARGET(HPMCOUNTER17)   \
`TARGET(HPMCOUNTER18)   \
`TARGET(HPMCOUNTER19)   \
`TARGET(HPMCOUNTER20)   \
`TARGET(HPMCOUNTER21)   \
`TARGET(HPMCOUNTER22)   \
`TARGET(HPMCOUNTER23)   \
`TARGET(HPMCOUNTER24)   \
`TARGET(HPMCOUNTER25)   \
`TARGET(HPMCOUNTER26)   \
`TARGET(HPMCOUNTER27)   \
`TARGET(HPMCOUNTER28)   \
`TARGET(HPMCOUNTER29)   \
`TARGET(HPMCOUNTER30)   \
`TARGET(HPMCOUNTER31)   \
`TARGET(HPMCOUNTER3H)   \
`TARGET(HPMCOUNTER4H)   \
`TARGET(HPMCOUNTER5H)   \
`TARGET(HPMCOUNTER6H)   \
`TARGET(HPMCOUNTER7H)   \
`TARGET(HPMCOUNTER8H)   \
`TARGET(HPMCOUNTER9H)   \
`TARGET(HPMCOUNTER10H)  \
`TARGET(HPMCOUNTER11H)  \
`TARGET(HPMCOUNTER12H)  \
`TARGET(HPMCOUNTER13H)  \
`TARGET(HPMCOUNTER14H)  \
`TARGET(HPMCOUNTER15H)  \
`TARGET(HPMCOUNTER16H)  \
`TARGET(HPMCOUNTER17H)  \
`TARGET(HPMCOUNTER18H)  \
`TARGET(HPMCOUNTER19H)  \
`TARGET(HPMCOUNTER20H)  \
`TARGET(HPMCOUNTER21H)  \
`TARGET(HPMCOUNTER22H)  \
`TARGET(HPMCOUNTER23H)  \
`TARGET(HPMCOUNTER24H)  \
`TARGET(HPMCOUNTER25H)  \
`TARGET(HPMCOUNTER26H)  \
`TARGET(HPMCOUNTER27H)  \
`TARGET(HPMCOUNTER28H)  \
`TARGET(HPMCOUNTER29H)  \
`TARGET(HPMCOUNTER30H)  \
`TARGET(HPMCOUNTER31H)  \
`TARGET(MVENDORID)      \
`TARGET(MARCHID)        \
`TARGET(MIMPID)         \
`TARGET(MHARTID)        \
`TARGET(MCONFIGPTR)     \
`TARGET(MSTATUS)        \
`TARGET(MSTATUSH)       \
`TARGET(MISA)           \
`TARGET(MIE)            \
`TARGET(MTVEC)          \
`TARGET(MSCRATCH)       \
`TARGET(MEPC)           \
`TARGET(MCAUSE)         \
`TARGET(MTVAL)          \
`TARGET(MIP)            \
`TARGET(MCYCLE)         \
`TARGET(MCYCLEH)        \
`TARGET(MINSTRET)       \
`TARGET(MINSTRETH)      \
`TARGET(MHPMCOUNTER3)   \
`TARGET(MHPMCOUNTER4)   \
`TARGET(MHPMCOUNTER5)   \
`TARGET(MHPMCOUNTER6)   \
`TARGET(MHPMCOUNTER7)   \
`TARGET(MHPMCOUNTER8)   \
`TARGET(MHPMCOUNTER9)   \
`TARGET(MHPMCOUNTER10)  \
`TARGET(MHPMCOUNTER11)  \
`TARGET(MHPMCOUNTER12)  \
`TARGET(MHPMCOUNTER13)  \
`TARGET(MHPMCOUNTER14)  \
`TARGET(MHPMCOUNTER15)  \
`TARGET(MHPMCOUNTER16)  \
`TARGET(MHPMCOUNTER17)  \
`TARGET(MHPMCOUNTER18)  \
`TARGET(MHPMCOUNTER19)  \
`TARGET(MHPMCOUNTER20)  \
`TARGET(MHPMCOUNTER21)  \
`TARGET(MHPMCOUNTER22)  \
`TARGET(MHPMCOUNTER23)  \
`TARGET(MHPMCOUNTER24)  \
`TARGET(MHPMCOUNTER25)  \
`TARGET(MHPMCOUNTER26)  \
`TARGET(MHPMCOUNTER27)  \
`TARGET(MHPMCOUNTER28)  \
`TARGET(MHPMCOUNTER29)  \
`TARGET(MHPMCOUNTER30)  \
`TARGET(MHPMCOUNTER31)  \
`TARGET(MHPMCOUNTER3H)  \
`TARGET(MHPMCOUNTER4H)  \
`TARGET(MHPMCOUNTER5H)  \
`TARGET(MHPMCOUNTER6H)  \
`TARGET(MHPMCOUNTER7H)  \
`TARGET(MHPMCOUNTER8H)  \
`TARGET(MHPMCOUNTER9H)  \
`TARGET(MHPMCOUNTER10H) \
`TARGET(MHPMCOUNTER11H) \
`TARGET(MHPMCOUNTER12H) \
`TARGET(MHPMCOUNTER13H) \
`TARGET(MHPMCOUNTER14H) \
`TARGET(MHPMCOUNTER15H) \
`TARGET(MHPMCOUNTER16H) \
`TARGET(MHPMCOUNTER17H) \
`TARGET(MHPMCOUNTER18H) \
`TARGET(MHPMCOUNTER19H) \
`TARGET(MHPMCOUNTER20H) \
`TARGET(MHPMCOUNTER21H) \
`TARGET(MHPMCOUNTER22H) \
`TARGET(MHPMCOUNTER23H) \
`TARGET(MHPMCOUNTER24H) \
`TARGET(MHPMCOUNTER25H) \
`TARGET(MHPMCOUNTER26H) \
`TARGET(MHPMCOUNTER27H) \
`TARGET(MHPMCOUNTER28H) \
`TARGET(MHPMCOUNTER29H) \
`TARGET(MHPMCOUNTER30H) \
`TARGET(MHPMCOUNTER31H) \
`TARGET(MCOUNTINHIBIT)  \
`TARGET(MHPMEVENT3)     \
`TARGET(MHPMEVENT4)     \
`TARGET(MHPMEVENT5)     \
`TARGET(MHPMEVENT6)     \
`TARGET(MHPMEVENT7)     \
`TARGET(MHPMEVENT8)     \
`TARGET(MHPMEVENT9)     \
`TARGET(MHPMEVENT10)    \
`TARGET(MHPMEVENT11)    \
`TARGET(MHPMEVENT12)    \
`TARGET(MHPMEVENT13)    \
`TARGET(MHPMEVENT14)    \
`TARGET(MHPMEVENT15)    \
`TARGET(MHPMEVENT16)    \
`TARGET(MHPMEVENT17)    \
`TARGET(MHPMEVENT18)    \
`TARGET(MHPMEVENT19)    \
`TARGET(MHPMEVENT20)    \
`TARGET(MHPMEVENT21)    \
`TARGET(MHPMEVENT22)    \
`TARGET(MHPMEVENT23)    \
`TARGET(MHPMEVENT24)    \
`TARGET(MHPMEVENT25)    \
`TARGET(MHPMEVENT26)    \
`TARGET(MHPMEVENT27)    \
`TARGET(MHPMEVENT28)    \
`TARGET(MHPMEVENT29)    \
`TARGET(MHPMEVENT30)    \
`TARGET(MHPMEVENT31)    \

`define CSRGEN__GENERATE_INTERFACE(csr) \
reg  [`ISA__XLEN-1:0] ``csr``_reg;   \
tri0 [`ISA__XLEN-1:0] ``csr``_in;    \
tri0                  ``csr``_write; \

`define CSRGEN__GENERATE_READ_ASSIGN(csr) \
assign reg_out = address == `CSR__``csr`` ? csr_interface.``csr``_reg : {`ISA__XLEN{1'bz}}; \
assign hit = address == `CSR__``csr`` ? 1'b1 : 1'bz;                                        \

`define CSRGEN__GENERATE_INITIAL_VALUE(csr) \
csr_interface.``csr``_reg <= `CSR__``csr``_VALUE; \

`define CSRGEN__GENERATE_WRITE(csr) \
if (csr_interface.``csr``_write) begin                                                                             \
    csr_interface.``csr``_reg <= csr_interface.``csr``_in;                                                         \
end else if (address == `CSR__``csr`` && write_reg) begin                                                          \
    csr_interface.``csr``_reg <= (value & `CSR__``csr``_MASK) | (csr_interface.``csr``_reg & ~`CSR__``csr``_MASK); \
end                                                                                                                \

`endif
